Universidad Tecnologica de El Salvador
Technological University of El Salvador
